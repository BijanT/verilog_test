module top (
    input i_sw,
    output o_led
    );

    thruwire tr(i_sw, o_led);

endmodule
